module signextend(b, a);

input [15:0] a;
output [31:0] b;

and Gate0(b[0],a[0],1);
and Gate1(b[1],a[1],1);
and Gate2(b[2],a[2],1);
and Gate3(b[3],a[3],1);
and Gate4(b[4],a[4],1);
and Gate5(b[5],a[5],1);
and Gate6(b[6],a[6],1);
and Gate7(b[7],a[7],1);
and Gate8(b[8],a[8],1);
and Gate9(b[9],a[9],1);
and Gate10(b[10],a[10],1);
and Gate11(b[11],a[11],1);
and Gate12(b[12],a[12],1);
and Gate13(b[13],a[13],1);
and Gate14(b[14],a[14],1);
and Gate15(b[15],a[15],1);
and Gate16(b[16],a[15],1);
and Gate17(b[17],a[15],1);
and Gate18(b[18],a[15],1);
and Gate19(b[19],a[15],1);
and Gate20(b[20],a[15],1);
and Gate21(b[21],a[15],1);
and Gate22(b[22],a[15],1);
and Gate23(b[23],a[15],1);
and Gate24(b[24],a[15],1);
and Gate25(b[25],a[15],1);
and Gate26(b[26],a[15],1);
and Gate27(b[27],a[15],1);
and Gate28(b[28],a[15],1);
and Gate29(b[29],a[15],1);
and Gate30(b[30],a[15],1);
and Gate31(b[31],a[15],1);


endmodule
