module bit32_2x1mux(A,B,S,ww);

input [31:0] A,B;
input S;

output [31:0] ww;



Two_One_Mux mux1(A[0],B[0],S,ww[0]);
Two_One_Mux mux2(A[1],B[1],S,ww[1]);
Two_One_Mux mux3(A[2],B[2],S,ww[2]);
Two_One_Mux mux4(A[3],B[3],S,ww[3]);
Two_One_Mux mux5(A[4],B[4],S,ww[4]);
Two_One_Mux mux6(A[5],B[5],S,ww[5]);
Two_One_Mux mux7(A[6],B[6],S,ww[6]);
Two_One_Mux mux8(A[7],B[7],S,ww[7]);
Two_One_Mux mux9(A[8],B[8],S,ww[8]);
Two_One_Mux mux10(A[9],B[9],S,ww[9]);
Two_One_Mux mux11(A[10],B[10],S,ww[10]);
Two_One_Mux mux12(A[11],B[11],S,ww[11]);
Two_One_Mux mux13(A[12],B[12],S,ww[12]);
Two_One_Mux mux14(A[13],B[13],S,ww[13]);
Two_One_Mux mux15(A[14],B[14],S,ww[14]);
Two_One_Mux mux16(A[15],B[15],S,ww[15]);
Two_One_Mux mux17(A[16],B[16],S,ww[16]);
Two_One_Mux mux18(A[17],B[17],S,ww[17]);
Two_One_Mux mux19(A[18],B[18],S,ww[18]);
Two_One_Mux mux20(A[19],B[19],S,ww[19]);
Two_One_Mux mux21(A[20],B[20],S,ww[20]);
Two_One_Mux mux22(A[21],B[21],S,ww[21]);
Two_One_Mux mux23(A[22],B[22],S,ww[22]);
Two_One_Mux mux24(A[23],B[23],S,ww[23]);
Two_One_Mux mux25(A[24],B[24],S,ww[24]);
Two_One_Mux mux26(A[25],B[25],S,ww[25]);
Two_One_Mux mux27(A[26],B[26],S,ww[26]);
Two_One_Mux mux28(A[27],B[27],S,ww[27]);
Two_One_Mux mux29(A[28],B[28],S,ww[28]);
Two_One_Mux mux30(A[29],B[29],S,ww[29]);
Two_One_Mux mux31(A[30],B[30],S,ww[30]);
Two_One_Mux mux32(A[31],B[31],S,ww[31]);





endmodule
