module sltModule(B,Output);

input B;
output [31:0] Output;

and Gate1(Output[0],1,B);
and Gate2(Output[1],0,0);
and Gate3(Output[2],0,0);
and Gate4(Output[3],0,0);
and Gate5(Output[4],0,0);
and Gate6(Output[5],0,0);
and Gate7(Output[6],0,0);
and Gate8(Output[7],0,0);
and Gate9(Output[8],0,0);
and Gate10(Output[9],0,0);
and Gate11(Output[10],0,0);
and Gate(Output[11],0,0);
and Gate12(Output[12],0,0);
and Gate13(Output[13],0,0);
and Gate14(Output[14],0,0);
and Gate15(Output[15],0,0);
and Gate16(Output[16],0,0);
and Gate17(Output[17],0,0);
and Gate18(Output[18],0,0);
and Gate19(Output[19],0,0);
and Gate20(Output[20],0,0);
and Gate21(Output[21],0,0);
and Gate22(Output[22],0,0);
and Gate23(Output[23],0,0);
and Gate24(Output[24],0,0);
and Gate25(Output[25],0,0);
and Gate26(Output[26],0,0);
and Gate27(Output[27],0,0);
and Gate28(Output[28],0,0);
and Gate29(Output[29],0,0);
and Gate30(Output[30],0,0);
and Gate31(Output[31],0,0);
	
endmodule
